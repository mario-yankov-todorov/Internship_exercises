module adder_with_feedback
     (
        // ------------------------------------------------------------------------------ 
        // Inputs and output 
        input    [16    -1:0]    in        ,
        output   [16    -1:0]    out       ,
        input                    reset     , 
        input                    clock   
        // ------------------------------------------------------------------------------
     );
		  
endmodule